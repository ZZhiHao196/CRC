// 自动生成的CRC配置文件
// 配置类型: mixed_two

`define CRC_WIDTH 'd8
`define CRC_POLY 'h17f
`define CRC_INIT 'hff
`define CRC_REFIN 'd0
`define CRC_REFOUT 'd1
`define CRC_XOROUT 'h0
