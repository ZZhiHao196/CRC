// 自动生成的CRC配置文件
// 配置类型: reflect

`define CRC_WIDTH 'd32
`define CRC_POLY 'h1d95f0ba3
`define CRC_INIT 'hffffffff
`define CRC_REFIN 'd1
`define CRC_REFOUT 'd1
`define CRC_XOROUT 'h0
