// 自动生成的CRC配置文件
// 配置类型: mixed_one

`define CRC_WIDTH 'd32
`define CRC_POLY 'h14d96321f
`define CRC_INIT 'hffffffff
`define CRC_REFIN 'd1
`define CRC_REFOUT 'd0
`define CRC_XOROUT 'h0
