// 自动生成的CRC配置文件
// 配置类型: standard

`define CRC_WIDTH 'd32
`define CRC_POLY 'h1e207f383
`define CRC_INIT 'hffffffff
`define CRC_REFIN 'd0
`define CRC_REFOUT 'd0
`define CRC_XOROUT 'h0
